module pisca (
		input clk,
		output led,
		input pow
);
